library verilog;
use verilog.vl_types.all;
entity alu_32_bit_vlg_vec_tst is
end alu_32_bit_vlg_vec_tst;
