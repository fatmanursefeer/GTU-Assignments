module not_32_bit (input [31:0] In, output [31:0] Out);

not not0 (Out[0], In[0]);
not not1 (Out[1], In[1]);
not not2 (Out[2], In[2]);
not not3 (Out[3], In[3]);
not not4 (Out[4], In[4]);
not not5 (Out[5], In[5]);
not not6 (Out[6], In[6]);
not not7 (Out[7], In[7]);
not not8 (Out[8], In[8]);
not not9 (Out[9], In[9]);
not not10 (Out[10], In[10]);
not not11 (Out[11], In[11]);
not not12 (Out[12], In[12]);
not not13 (Out[13], In[13]);
not not14 (Out[14], In[14]);
not not15 (Out[15], In[15]);
not not16 (Out[16], In[16]);
not not17 (Out[17], In[17]);
not not18 (Out[18], In[18]);
not not19 (Out[19], In[19]);
not not20 (Out[20], In[20]);
not not21 (Out[21], In[21]);
not not22 (Out[22], In[22]);
not not23 (Out[23], In[23]);
not not24 (Out[24], In[24]);
not not25 (Out[25], In[25]);
not not26 (Out[26], In[26]);
not not27 (Out[27], In[27]);
not not28 (Out[28], In[28]);
not not29 (Out[29], In[29]);
not not30 (Out[30], In[30]);
not not31 (Out[31], In[31]);

endmodule
